library IEEE;
use IEEE.std_logic_1164.all;  
use IEEE.numeric_std.all;     
use IEEE.std_logic_textio.all; 
library STD;    
use STD.textio.all;

library psx;

entity etb  is
end entity;

architecture arch of etb is

   signal clk1x               : std_logic := '1';
   signal clk2x               : std_logic := '1';
            
   signal reset               : std_logic := '1';
   
   signal clk1xToggle         : std_logic := '0';
   signal clk1xToggle2X       : std_logic := '0';
   signal clk2xIndex          : std_logic := '0';
   
   -- gte
   signal gte_busy            : std_logic;
   signal gte_readAddr        : unsigned(5 downto 0) := (others => '0');
   signal gte_readData        : unsigned(31 downto 0);
   signal gte_writeAddr       : unsigned(5 downto 0);
   signal gte_writeData       : unsigned(31 downto 0);
   signal gte_writeEna        : std_logic; 
   signal gte_cmdData         : unsigned(31 downto 0);
   signal gte_cmdEna          : std_logic; 
   
   -- testbench
   signal cmdCount            : integer := 0;
   
begin

   clk1x  <= not clk1x  after 15 ns;
   clk2x  <= not clk2x  after 7500 ps;
   
   reset  <= '0' after 3000 ns;
   
   -- clock index
   process (clk1x)
   begin
      if rising_edge(clk1x) then
         clk1xToggle <= not clk1xToggle;
      end if;
   end process;
   
   process (clk2x)
   begin
      if rising_edge(clk2x) then
         clk1xToggle2x <= clk1xToggle;
         clk2xIndex    <= '0';
         if (clk1xToggle2x = clk1xToggle) then
            clk2xIndex <= '1';
         end if;
      end if;
   end process;
   
   igte : entity psx.gte
   port map
   (
      clk2x                => clk2x,     
      clk2xIndex           => clk2xIndex,
      ce                   => '1',        
      reset                => reset,     
      
      gte_busy             => gte_busy,     
      gte_readAddr         => gte_readAddr, 
      gte_readData         => gte_readData, 
      gte_writeAddr        => gte_writeAddr,
      gte_writeData        => gte_writeData,
      gte_writeEna         => gte_writeEna, 
      gte_cmdData          => gte_cmdData,  
      gte_cmdEna           => gte_cmdEna  
   );
   
   process
      file infile          : text;
      variable f_status    : FILE_OPEN_STATUS;
      variable inLine      : LINE;
      variable para_type   : std_logic_vector(7 downto 0);
      variable para_addr   : std_logic_vector(7 downto 0);
      variable para_data   : std_logic_vector(31 downto 0);
      variable space       : character;
   begin
      
      gte_writeEna <= '0';
      gte_cmdEna   <= '0';
      
      wait until reset = '0';
         
      file_open(f_status, infile, "R:\gte_test_fpsxa.txt", read_mode);
      
      while (not endfile(infile)) loop
         
         readline(infile,inLine);
         
         HREAD(inLine, para_type);
         Read(inLine, space);
         HREAD(inLine, para_addr);
         Read(inLine, space);
         HREAD(inLine, para_data);
         
         if (para_type = x"01") then
            gte_cmdData <= unsigned(para_data);
            gte_cmdEna  <= '1';
         elsif (para_type = x"02") then
            gte_writeAddr <= unsigned(para_addr(5 downto 0));
            gte_writeData <= unsigned(para_data);
            gte_writeEna  <= '1';
         end if;
         
         cmdCount <= cmdCount + 1;
         wait until rising_edge(clk1x);
         
         gte_writeEna <= '0';
         gte_cmdEna   <= '0';
         
         while (gte_busy = '1') loop
            wait until rising_edge(clk1x);
         end loop;
         
      end loop;
      
      file_close(infile);
      
      wait for 1 us;
      
      if (cmdCount >= 0) then
         report "DONE" severity failure;
      end if;
      
      
   end process;
   
   
end architecture;


